`timescale 1ns / 1ps

module Bus_mux(
input [1:0] bus_grant,
input [1:0] slave_sel 
    );
endmodule
